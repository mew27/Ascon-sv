module ascon_ps (
  ports
);
  
endmodule
