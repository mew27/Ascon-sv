module ascon;
`timescale 1ns/1ps

initial begin
  $display("Hello World in System Verilog!");
  #10;
  $finish;
end  

endmodule
